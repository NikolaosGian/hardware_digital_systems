`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:47:47 12/05/2021 
// Design Name: 
// Module Name:    dec5to32 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dec5to32(
    input [4:0] enc,
    output reg [31:0] dec
    );

always @(*) begin

case (enc)
	
	5'b00000: dec = 32'h0000_0001;
	5'b00001: dec = 32'h0000_0002;
	5'b00010: dec = 32'h0000_0004;
	5'b00011: dec = 32'h0000_0008;
	5'b00100: dec = 32'h0000_0010;
	5'b00101: dec = 32'h0000_0020;
	5'b00110: dec = 32'h0000_0040;
	5'b00111: dec = 32'h0000_0080;
	5'b01000: dec = 32'h0000_0100;
	5'b01001: dec = 32'h0000_0200;
	5'b01010: dec = 32'h0000_0400;
	5'b01011: dec = 32'h0000_0800;
	5'b01100: dec = 32'h0000_1000;
	5'b01101: dec = 32'h0000_2000;
	5'b01110: dec = 32'h0000_4000;
	5'b01111: dec = 32'h0000_8000;
	5'b10000: dec = 32'h0001_0000;
	5'b10001: dec = 32'h0002_0000;
	5'b10010: dec = 32'h0004_0000;
	5'b10011: dec = 32'h0008_0000;
	5'b10100: dec = 32'h0010_0000;
	5'b10101: dec = 32'h0020_0000;
	5'b10110: dec = 32'h0040_0000;
	5'b10111: dec = 32'h0080_0000;
	5'b11000: dec = 32'h0100_0000;
	5'b11001: dec = 32'h0200_0000;
	5'b11010: dec = 32'h0400_0000;
	5'b11011: dec = 32'h0800_0000;
	5'b11100: dec = 32'h1000_0000;
	5'b11101: dec = 32'h2000_0000;
	5'b11110: dec = 32'h4000_0000;
	5'b11111: dec = 32'h8000_0000;
	
endcase

end

endmodule
